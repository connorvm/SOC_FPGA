This file will be handling the status resgiter logic