-- This file will handle all of the opcodes and its operations

-- Authors: Connor Van Meter, Alex Salois


    library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    use IEEE.NUMERIC_STD.ALL;
    use IEEE.std_logic_unsigned.all;
    
    LIBRARY altera;
    USE altera.altera_primitives_components.all;
    
    
    entity operations is
        port(
            clk            : in  std_logic;                         -- system clock
            reset          : in  std_logic;                         -- system reset
            PB             : in  std_logic;                         -- Pushbutton to change state  
            SW             : in  std_logic_vector(3 downto 0);      -- Switches that determine next state
            HS_LED_control : in  std_logic;                         -- Software is in control when asserted (=1)
            SYS_CLKs_sec   : in  std_logic_vector(31 downto 0);     -- Number of system clock cycles in one second
            Base_rate      : in  std_logic_vector(7 downto 0);      -- base transition time in seconds, fixed-point data type
            LED_reg        : in  std_logic_vector(7 downto 0);      -- LED register
            LED            : out std_logic_vector(7 downto 0)       -- LEDs on the DE10-Nano board
        );
    end entity operations;
    
    
    architecture operations_arch of operations is


        begin



    end architecture operations_arch;
    