This file will be the top level in our design
