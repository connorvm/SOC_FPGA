Make this work

