This file will handle all of the opcodes and its operations