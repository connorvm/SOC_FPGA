-- Authors: Connor Van Meter & Alex Salois
-- EELE 468

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;

entity add_1 is
  port (Input  : in  std_logic_vector (7 downto 0);
	Output : out std_logic_vector (7 downto 0));
end entity;

architecture add_1_arch of add_1 is

  begin



end architecture;